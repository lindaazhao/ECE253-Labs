module part3(A, B, Function, ALUout);
endmodule